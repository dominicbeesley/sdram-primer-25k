-- MIT License
-- -----------------------------------------------------------------------------
-- Copyright (c) 2024 Dominic Beesley https://github.com/dominicbeesley
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
-- ----------------------------------------------------------------------

-- Company: 			Dossytronics
-- Engineer: 			Dominic Beesley
-- 
-- Create Date:    	22/05/2024
-- Design Name: 
-- Module Name:    	fb_port_io
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 		fishbone bus - a simple 8 bit input/output port
-- Dependencies: 
--
-- Revision: 
-- Additional Comments: 
--
----------------------------------------------------------------------------------



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

library work;
use work.fishbone.all;
use work.common.all;

entity fb_port_io is
	generic (
		SIM								: boolean := false;							-- skip some stuff, i.e. slow sdram start up
		CLOCKSPEED						: natural										-- fast clock speed in mhz						
	);
	port(

		-- fishbone signals
		fb_syscon_i						: in 	fb_syscon_t;
		fb_c2p_i							: in 	fb_con_o_per_i_t;
		fb_p2c_o							: out fb_con_i_per_o_t;

		-- serial
		bits_o							: out std_logic_vector(7 downto 0);
		bits_i							: in  std_logic_vector(7 downto 0)
	);
end fb_port_io;

architecture rtl of fb_port_io is
	
begin

	fb_p2c_o.rdy <= '1';
	fb_p2c_o.stall <= '0';
	fb_p2c_o.D_rd <= bits_i;

	p_fb:process(fb_syscon_i)
	variable v_we : std_logic;
	variable v_cyc: std_logic;
	begin
		if fb_syscon_i.rst = '1' then
			bits_o <= (others => '0');
			v_we := '0';
			v_cyc := '0';
		elsif rising_edge(fb_syscon_i.clk) then
			if fb_c2p_i.cyc = '1' and fb_c2p_i.a_stb = '1' then
				v_cyc := '1';
				v_we := fb_c2p_i.we;
			end if;

			if v_cyc then
				if v_we = '0' then
					fb_p2c_o.ack <= '1';
					v_cyc := '0';
				elsif v_we = '1' and fb_c2p_i.d_wr_stb = '1' then
					fb_p2c_o.ack <= '1';
					bits_o <= fb_c2p_i.d_wr;
					v_cyc := '0';
				end if;
			end if;
		end if;
	end process;

end rtl;